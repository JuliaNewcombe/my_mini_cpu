module not_val (input [31:0] A, output [31:0] result);
	
	assign result = ~A;
	
endmodule